
package complex_pkg;

	localparam logic [ 0:0 ]
		RE = 0,
		IM = 1;

endpackage: complex_pkg

