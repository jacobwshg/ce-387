
module background_sub(

);

endmodule

