
module fft_stage #(
	IDX_WIDTH = 5,
	IDX_SIZE  = 2 ** IDX_WIDTH,
	DATA_WIDTH = 32
)
(
	
);

endmodule: fft_stage

