
module matmul_tb();

endmodule

