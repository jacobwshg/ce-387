
module highlight(

);

endmodule

