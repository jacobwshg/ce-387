
module grayscale(

);

endmodule

